module models
