module models

pub const allowed_post_type = ['post', 'page']

pub const allowed_post_status = ['published', 'draft', 'scheduled']

pub const allowed_visibility = ['public', 'paid']

pub const allowed_role = ['admin', 'member', 'developer', 'author', 'contributor']
