module models

pub const allowed_post_status = ['published', 'draft', 'scheduled']

pub const allowed_visibility = ['public', 'paid']
