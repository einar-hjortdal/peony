module models

// customer.id can be taken with SELECT BIN_TO_UUID("id", 0)
// customer.id can be stored as UUID_TO_BIN(, 0)
