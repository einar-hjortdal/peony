module redis
// TODO implement bullmq-like queue

// fn create new queue with given name
// method add item (json string) to named queue
// create concurrent worker
// listen to events: job completions