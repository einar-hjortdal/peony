module redis
// TODO implement event bus